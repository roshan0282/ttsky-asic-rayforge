module asic(

);


endmodule