/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_asic (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  wire rst;
  wire [9:0] clk_per_bit;

  assign clk_per_bit = {uio_in[7:0], 2'b00}; // set upper 8 bits
  assign rst = ~rst_n;
  assign uio_oe = 8'b0000_0000; // set bidirectional as inputs
  assign uio_out = 8'b0000_0000; // set unused bidirectional outputs to LOW

  asic asic0(.in(ui_in),.out(uo_out));
  // List all unused inputs to prevent warnings
  wire _unused = &{ui_in[7:1], ena, 1'b0};

endmodule
